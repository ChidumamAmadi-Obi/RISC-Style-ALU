`include "ALU_constants.svh"

`timescale 1ns/1ps // specifies the time units and precision for sim

module test;

endmodule
